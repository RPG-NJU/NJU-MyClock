module AlarmRun(
	);
	
endmodule
